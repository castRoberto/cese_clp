library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

--=============================================================================

entity fir is

  generic (
	  C_DATA_W  : natural := 12
	);

  port (
    clk     : in std_logic;
    fsclk   : in std_logic;
    rst     : in std_logic;
    x_in    : in unsigned (C_DATA_W - 1 downto 0);
    y_out   : out unsigned (C_DATA_W * 2 - 1 downto 0)
  );

end fir;

--=============================================================================

architecture fir_arc of fir is

  constant C_TAPS : natural := 51;  -- número de coeficientes

  type state_machine is (idle_st, active_st);

  type t_data_array is array (0 to C_TAPS - 1)
                     of signed (C_DATA_W - 1 downto 0);

  signal delay_line : t_data_array := (others => (others => '0'));

  signal coeffs : t_data_array := (
    to_signed( 105, C_DATA_W),
    to_signed(  74, C_DATA_W),
    to_signed(-112, C_DATA_W),
    to_signed( -53, C_DATA_W),
    to_signed(  -5, C_DATA_W),
    to_signed( -76, C_DATA_W),
    to_signed(   2, C_DATA_W),
    to_signed( -30, C_DATA_W),
    to_signed( -40, C_DATA_W),
    to_signed(  22, C_DATA_W),
    to_signed( -54, C_DATA_W),
    to_signed(  10, C_DATA_W),
    to_signed(   0, C_DATA_W),
    to_signed( -50, C_DATA_W),
    to_signed(  51, C_DATA_W),
    to_signed( -52, C_DATA_W),
    to_signed(   3, C_DATA_W),
    to_signed(  41, C_DATA_W),
    to_signed( -92, C_DATA_W),
    to_signed(  94, C_DATA_W),
    to_signed( -54, C_DATA_W),
    to_signed( -50, C_DATA_W),
    to_signed( 181, C_DATA_W),
    to_signed(-324, C_DATA_W),
    to_signed( 423, C_DATA_W),
    to_signed(1583, C_DATA_W),
    to_signed( 423, C_DATA_W),
    to_signed(-324, C_DATA_W),
    to_signed( 181, C_DATA_W),
    to_signed( -50, C_DATA_W),
    to_signed( -54, C_DATA_W),
    to_signed(  94, C_DATA_W),
    to_signed( -92, C_DATA_W),
    to_signed(  41, C_DATA_W),
    to_signed(   3, C_DATA_W),
    to_signed( -52, C_DATA_W),
    to_signed(  51, C_DATA_W),
    to_signed( -50, C_DATA_W),
    to_signed(   0, C_DATA_W),
    to_signed(  10, C_DATA_W),
    to_signed( -54, C_DATA_W),
    to_signed(  22, C_DATA_W),
    to_signed( -40, C_DATA_W),
    to_signed( -30, C_DATA_W),
    to_signed(   2, C_DATA_W),
    to_signed( -76, C_DATA_W),
    to_signed(  -5, C_DATA_W),
    to_signed( -53, C_DATA_W),
    to_signed(-112, C_DATA_W),
    to_signed(  74, C_DATA_W),
    to_signed( 105, C_DATA_W)
  );

  signal state : state_machine := idle_st;

  signal counter : integer range 0 to C_TAPS - 1 := C_TAPS - 1;

  signal output : signed (C_DATA_W * 2 - 1 downto 0) := (others=>'0');

  signal accumulator : signed (C_DATA_W * 2 - 1 downto 0) := (others=>'0');

  signal fsclk_q : std_logic := '0';

begin

  --
  y_out <= unsigned (std_logic_vector(output));

  --
  fir : process (clk)

    variable sum_v : signed (C_DATA_W * 2 - 1 downto 0) := (others=>'0');

  begin

    if rising_edge(clk) then

      fsclk_q <= fsclk;

      case state is

        when idle_st =>

          if fsclk = '1' and fsclk_q = '0' then

            state <= active_st;

          end if;

        when active_st =>

          if counter > 0 then

            counter <= counter - 1;

          else

            counter <= C_TAPS - 1;
            state <= idle_st;

          end if;

          -- Shifting the delay line
          --
          if counter > 0 then

            delay_line (counter) <= delay_line (counter - 1);

          else

            delay_line (counter) <= signed (std_logic_vector (x_in));

          end if;

          -- Multiplying the delay line with coefficients
          --
          if counter > 0 then

            sum_v := delay_line (counter) * coeffs (counter);
            accumulator <= accumulator + sum_v;

          else

            accumulator <= (others=>'0');
            sum_v := delay_line (counter) * coeffs (counter);
            output <= accumulator + sum_v;

          end if;

      end case;

    end if;

  end process;

end;

--=============================================================================